** Profile: "SCHEMATIC1-sim1"  [ i:\ee\semester_2\circuits\lab\ec_report-main\report 5\pspice\sim-schematic1-sim1.sim ] 

** Creating circuit file "sim-schematic1-sim1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V2 -100 100 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\sim-SCHEMATIC1.net" 


.END
