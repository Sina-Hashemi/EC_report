** Profile: "SCHEMATIC1-sim"  [ I:\EE\semester_2\circuits\Lab\EC_report-main\Report 3\Pspice\pspice-SCHEMATIC1-sim.sim ] 

** Creating circuit file "pspice-SCHEMATIC1-sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of E:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 1 10000
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pspice-SCHEMATIC1.net" 


.END
